//*****************************************************
// Project		: Assignment 1
// File			: section2_a1
// Editor		: Wenmei Wang
// Date			: 15/10/2024
// Description	: Assignment 1
//*****************************************************

module ha (

	input	a, b,
	output	s, c
	
);

	assign s = a ^ b;
	assign c = a & b;

endmodule